wire clk  = i_gen_external_clk_0.clk;
wire rstnn = i_gen_external_clk_0.rstnn;
wire external_rstnn = rstnn;
