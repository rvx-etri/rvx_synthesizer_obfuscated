`include "user_ddr3_body.vh"
