`include "ervp_global.vh"
`include "ervp_endian.vh"
`include "ervp_axi_define.vh"
`include "ervp_ahb_define.vh"

`include "ervp_platform_controller_memorymap_offset.vh"
`include "ervp_jtag_memorymap_offset.vh"
`include "ervp_mmiox1_memorymap_offset.vh"

`include "platform_info.vh"
`include "sim_info.vh"
`include "hex_size.vh"

`include "timescale.vh"
