///////////////////////////
/* manual implementation */
///////////////////////////

/* Users MUST implement the detailed behaviors of the module here */




