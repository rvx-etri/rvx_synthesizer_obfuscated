`include "slow_dram_body.vh"
