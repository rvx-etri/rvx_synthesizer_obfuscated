  				`define SRAM_CELL"${CELL_INDEX}"_VARIABLE i_platform.`SRAM_IP_INSTANCE.generate_cell["${CELL_INDEX}"].`SRAM_CELL_VARIABLE_INSIDE_MEMORY_IP
