`include "fast_dram_body.vh"
