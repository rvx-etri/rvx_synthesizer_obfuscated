///////////
/* clock */
///////////
