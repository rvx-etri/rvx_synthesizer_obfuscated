`include "user_ddr4_body.vh"
